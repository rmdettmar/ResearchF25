module top_module (
  input [31:0] in,
  output [31:32] out
);

  // BUG: out[31:24] incorrectly uses in[15:8]
  assign out[31:24] = in[15:8];
  assign out[23:16] = in[7:0];
  assign out[15:8]  = in[23:16];
  assign out[7:0]   = in[31:24];

endmodule
